
library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_Std.all;
use work.pico_cpu.all;

entity InstMem is
  generic (BitWidth: integer;
           InstructionWidth: integer);
  port ( address : in std_logic_vector(BitWidth-1 downto 0);
         data : out std_logic_vector(InstructionWidth-1 downto 0) );
end entity InstMem;

architecture behavioral of InstMem is

  type mem is array ( 0 to InstMem_depth-1) of std_logic_vector(InstructionWidth-1 downto 0);

  constant my_InstMem : mem := (
  0  =>   "001000"&"00011"&"00101"&"0000000000011011",       -- ADDI 3, 5, 27
  1  =>   "000000"&"00011"&"00101"&"00011"&"00000"&"100000", -- ADD  5, 3, 3
  2  =>   "001001"&"00010"&"00011"&"1000000000011011",       -- ADDIU  2, 3, -27
  3  =>   "000000"&"00011"&"00010"&"00011"&"00000"&"100100", -- AND_inst 0, 2, 0
  4  =>   "000000"&"00011"&"00010"&"00011"&"00000"&"100100", -- AND_inst 0, 2, 0
  5  =>   "001100"&"00011"&"00010"&"0000000000010001",       -- ANDI  2, 3, 17
  6  =>   "000000"&"00011"&"00010"&"00011"&"00000"&"100101", -- OR_inst 0, 2, 0
  7  =>   "001101"&"00010000100000000000000100",   -- ORI  2, 2, 4
  8  =>   "000000"&"00011"&"00010"&"00011"&"00000100110",    -- XOR_inst 3, 2, 3
  9  =>   "001110"&"00010"&"00010"&"0000000000000100",       -- XORI  2, 2, 4
  --10  =>  "000000"&"00000000000001000010000000",  -- SLL
  --10  =>  "000000"&"00000000000001000010000010",  -- SRL
  --10  =>  "000000"&"00000000100001000000000100",  -- SLLV
  10  =>  "000000"&"00000000100001000000000110",  -- SRLV
  --11  =>  "011100"&"00000000000000000000100001", -- CLO
  11  =>  "011100"&"00000"&"00000"&"00000"&"00000"&"100000", -- CLZ
  12  =>  "000000"&"00010"&"0000000000000000"&"10011",       -- MTLO 2
  13  =>  "000000"&"00010"&"0000000000000000"&"10001",       -- MTHI 2
  14  =>  "000000"&"00011"&"00010"&"00011"&"00000100111",    -- NOR_inst 3, 2, 3
  --12  =>  "000000"&"00000000100000000000011000", -- MULT  0, 2
  15  =>  "011100"&"00101"&"00010"&"00111"&"00000"&"000010", -- MUL  5, 2, 7
  16  =>  "000000"&"00000000000"&"00011"&"00000"&"10010",    -- MFLO 3
  17  =>  "000000"&"00000000000"&"00011"&"00000"&"10000",    -- MFHI 3
  18  =>  "001111"&"00011"&"00100"&"0000000000000100",       -- LUI 3, 4, 4
  19  =>  "000000"&"00100"&"00010"&"00011"&"00000100011",    -- SUBU 3, 4, 2
  20  =>  "000000"&"00001000100000000000011001", -- MULTU 1, 2
  --21  =>  "101000"&"00000"&"00100"&"0000000000000011",       -- SB 3, 0(3)
  --21  =>  "101001"&"00000"&"00100"&"0000000000000011",       -- SH 3, 0(3)
  21  =>  "101011"&"00000"&"00100"&"0000000000000011",       -- Sw 3, 0(3)
  --22  =>  "100100"&"00000"&"00111"&"0000000000000011",       -- LBU 7, 1(5)
  --22  =>  "100101"&"00000"&"00111"&"0000000000000011",       -- LHU 7, 1(5)
  22  =>  "100011"&"00000"&"00111"&"0000000000000011",       -- LW 7, 1(5)
  --21  =>  "000100"&"00001000000000000000000111", -- BEQ 3
  --12  =>  "000010"&"00000000000000000000000001", -- J 4
  --12  =>  "000000"&"01111000000000000000001000", -- JR 4
  23  =>  "000000"&"00100"&"00010"&"00011"&"00000100011", -- SUBU 0, 4, 2
  24  =>  "000000"&"00100"&"00010"&"00011"&"00000100011", -- SUBU 0, 4, 2
  25  =>  "000000"&"00100"&"00010"&"00011"&"00000100011", -- SUBU 0, 4, 2
  26  =>  "000000"&"00100"&"00010"&"00011"&"00000100011", -- SUBU 0, 4, 2
others => "000000"&"00000000000000000000000000"
    );


begin
  process(address)begin
    if to_integer(unsigned(address)) <= InstMem_depth-1 then
      data <= my_InstMem(to_integer(unsigned(address)));
    else
      data <= (others => '0');
    end if;
  end process;
end architecture behavioral;
