
library ieee;
use ieee.std_logic_1164.all;
use IEEE.Numeric_Std.all;
use work.pico_cpu.all;

entity InstMem is
  generic (BitWidth: integer;
           InstructionWidth: integer);
  port ( address : in std_logic_vector(BitWidth-1 downto 0);
         data : out std_logic_vector(InstructionWidth-1 downto 0) );
end entity InstMem;

architecture behavioral of InstMem is

  type mem is array ( 0 to InstMem_depth-1) of std_logic_vector(InstructionWidth-1 downto 0);

  constant my_InstMem : mem := (
0  =>   "10000100000000000000000000000000011000",--Load_R0_Dir   R0 = 24
1  =>   "00111100000000000000000000000000000000",--OR_A_R0       ACC = 24
2  =>   "00011000000000000000000000000000000000",--IncA         ACC = 25
3  =>   "00001100000000000000000000000000000000",--Sub_A_R0      ACC = 1
4  =>   "11111000000000000000000000000000000000",--NOP
5  =>   "01011000000000000000000000000000001001",--JmpC 7        Jump
6  =>   "11111000000000000000000000000000000000",--NOP
7  =>   "11111000000000000000000000000000000000",--NOP
8  =>   "11111000000000000000000000000000000000",--NOP
9  =>   "11111000000000000000000000000000000000",--NOP
10 =>   "00110000000000000000000000000000000000",--RRC
11 =>   "00110100000000000000000000000000000000",--RLC          ACC = 1
12 =>   "11111000000000000000000000000000000000",--NOP
13 =>   "01101100000000000000000000000000000000",--ClearC
14 =>   "10000000000000000000000000000000010000",--Store_A_Mem   MEM[16] = 1
15 =>   "11110000000000000000000000000000000000",--PUSH
16 =>   "01111000000000000000000000000000000000",--SavePC
17 =>   "11110000000000000000000000000000000000",--PUSH
18 =>   "01001100000000000000000000000000011010",--Jmp 23
19 =>   "11111000000000000000000000000000000000",--NOP
20 =>   "11111000000000000000000000000000000000",--NOP
21 =>   "11111000000000000000000000000000000000",--NOP
22 =>   "11110100000000000000000000000000000000", --pop
23 =>   "00100100000000000000000000000000000000", --ShiftArithL
24 =>   "00011100000000000000000000000000000000",--DecA
25 =>   "11111100000000000000000000000000000000", --HALT
26 =>   "01111100000000000000000000000000010000",--Load_A_Mem
27 =>   "00111000000000000000000000000000000000",--AND
28 =>   "01010000000000000000000000000000011011",--JMPZ 27
29 =>   "11111000000000000000000000000000000000",--NOP
30 =>   "01101100000000000000000000000000000000",--ClearZ
31 =>   "00000100000000000000000000000000010000",--Add_A_Mem
32 =>   "00010000000000000000000000000000010000",--Sub_A_Mem
33 =>   "00000000000000000000000000000000000000",--ADD_A_B
34 =>   "00010100000000000000000000000000001100",--SUB_A_DIR C
35 =>   "01000100000000000000000000000000000000",--FlipA
36 =>   "01000000000000000000000000000000000000",--XOR_A_B
37 =>   "01001000000000000000000000000000000000",--NegA
38 =>   "00100000000000000000000000000000000000",--ShiftArithR
39 =>   "00101100000000000000000000000000000000",--ShiftA_L
40 =>   "00101000000000000000000000000000000000",--ShiftA_R
41 =>   "01110000000000000000000000000000000000",--ClearACC
42 =>   "11110100000000000000000000000000000000",--POP
43 =>   "11111000000000000000000000000000000000",--NOP
44 =>   "11111000000000000000000000000000000000",--NOP
45 =>   "11111000000000000000000000000000000000",--NOP
46 =>   "00001000000000000000000000000000000110",--Add_A_Dir
47 =>   "11111000000000000000000000000000000000",--NOP
48 =>   "11111000000000000000000000000000000000",--NOP
49 =>   "01110100000000000000000000000000000000",--LoadPC
others => "00000000000000000000000000000000000000"
    );


begin
  process(address)begin
    if to_integer(unsigned(address)) <= InstMem_depth-1 then
      data <= my_InstMem(to_integer(unsigned(address)));
    else
      data <= (others => '0');
    end if;
  end process;
end architecture behavioral;
